<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-95.1665,15.25,222.467,-141.75</PageViewport>
<gate>
<ID>2</ID>
<type>BE_JKFF_LOW_NT</type>
<position>44,-26</position>
<input>
<ID>J</ID>9 </input>
<input>
<ID>K</ID>9 </input>
<output>
<ID>Q</ID>15 </output>
<input>
<ID>clock</ID>1 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4</ID>
<type>BB_CLOCK</type>
<position>26,-26</position>
<output>
<ID>CLK</ID>1 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>10</ID>
<type>BE_JKFF_LOW_NT</type>
<position>56,-26</position>
<input>
<ID>J</ID>11 </input>
<input>
<ID>K</ID>11 </input>
<output>
<ID>Q</ID>19 </output>
<input>
<ID>clock</ID>16 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>11</ID>
<type>BE_JKFF_LOW_NT</type>
<position>70,-26</position>
<input>
<ID>J</ID>6 </input>
<input>
<ID>K</ID>6 </input>
<output>
<ID>Q</ID>10 </output>
<input>
<ID>clock</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>12</ID>
<type>AA_TOGGLE</type>
<position>13.5,14</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>14</ID>
<type>DE_TO</type>
<position>24.5,14</position>
<input>
<ID>IN_0</ID>7 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 1</lparam></gate>
<gate>
<ID>16</ID>
<type>DA_FROM</type>
<position>33.5,-21.5</position>
<input>
<ID>IN_0</ID>9 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 1</lparam></gate>
<gate>
<ID>19</ID>
<type>DA_FROM</type>
<position>65,-21</position>
<input>
<ID>IN_0</ID>6 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID 1</lparam></gate>
<gate>
<ID>23</ID>
<type>GA_LED</type>
<position>60.5,-24</position>
<input>
<ID>N_in0</ID>19 </input>
<input>
<ID>N_in1</ID>18 </input>
<input>
<ID>N_in3</ID>13 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>25</ID>
<type>GA_LED</type>
<position>71.5,-21</position>
<input>
<ID>N_in0</ID>10 </input>
<input>
<ID>N_in3</ID>14 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>26</ID>
<type>DA_FROM</type>
<position>52,-21</position>
<input>
<ID>IN_0</ID>11 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID 1</lparam></gate>
<gate>
<ID>30</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>78.5,-13.5</position>
<input>
<ID>IN_0</ID>17 </input>
<input>
<ID>IN_1</ID>13 </input>
<input>
<ID>IN_2</ID>14 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 6</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>32</ID>
<type>GA_LED</type>
<position>49,-24</position>
<input>
<ID>N_in0</ID>15 </input>
<input>
<ID>N_in1</ID>16 </input>
<input>
<ID>N_in3</ID>17 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>34</ID>
<type>AA_LABEL</type>
<position>46,-4.5</position>
<gparam>LABEL_TEXT 1) ASYNC 3-bit up-counter using -ve edge triggered JK-FF</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>48</ID>
<type>AA_LABEL</type>
<position>46.5,-37</position>
<gparam>LABEL_TEXT 2) ASYNC 3-bit down-counter using -ve edge triggered JK-FF</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>72</ID>
<type>BB_CLOCK</type>
<position>21.5,-55</position>
<output>
<ID>CLK</ID>67 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>73</ID>
<type>BE_JKFF_LOW_NT</type>
<position>32,-55</position>
<input>
<ID>J</ID>68 </input>
<input>
<ID>K</ID>68 </input>
<output>
<ID>Q</ID>70 </output>
<input>
<ID>clock</ID>67 </input>
<output>
<ID>nQ</ID>73 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>74</ID>
<type>DA_FROM</type>
<position>26.5,-50</position>
<input>
<ID>IN_0</ID>68 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 1</lparam></gate>
<gate>
<ID>75</ID>
<type>DA_FROM</type>
<position>39.5,-49.5</position>
<input>
<ID>IN_0</ID>69 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 1</lparam></gate>
<gate>
<ID>76</ID>
<type>BE_JKFF_LOW_NT</type>
<position>45,-54.5</position>
<input>
<ID>J</ID>69 </input>
<input>
<ID>K</ID>69 </input>
<output>
<ID>Q</ID>71 </output>
<input>
<ID>clock</ID>73 </input>
<output>
<ID>nQ</ID>74 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>77</ID>
<type>DA_FROM</type>
<position>53,-49.5</position>
<input>
<ID>IN_0</ID>75 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 1</lparam></gate>
<gate>
<ID>78</ID>
<type>BE_JKFF_LOW_NT</type>
<position>58.5,-54.5</position>
<input>
<ID>J</ID>75 </input>
<input>
<ID>K</ID>75 </input>
<output>
<ID>Q</ID>72 </output>
<input>
<ID>clock</ID>74 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>79</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>68.5,-45.5</position>
<input>
<ID>IN_0</ID>70 </input>
<input>
<ID>IN_1</ID>71 </input>
<input>
<ID>IN_2</ID>72 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 6</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>81</ID>
<type>BB_CLOCK</type>
<position>18,-87.5</position>
<output>
<ID>CLK</ID>76 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>82</ID>
<type>BE_JKFF_LOW_NT</type>
<position>37.5,-87.5</position>
<input>
<ID>J</ID>77 </input>
<input>
<ID>K</ID>77 </input>
<output>
<ID>Q</ID>106 </output>
<input>
<ID>clock</ID>76 </input>
<output>
<ID>nQ</ID>86 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>83</ID>
<type>DA_FROM</type>
<position>19,-82.5</position>
<input>
<ID>IN_0</ID>77 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 1</lparam></gate>
<gate>
<ID>89</ID>
<type>AA_LABEL</type>
<position>47,-66</position>
<gparam>LABEL_TEXT 3) ASYNC 3-bit up/down-counter using -ve edge triggered JK-FF</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>91</ID>
<type>AA_AND2</type>
<position>48.5,-84.5</position>
<input>
<ID>IN_0</ID>100 </input>
<input>
<ID>IN_1</ID>106 </input>
<output>
<ID>OUT</ID>88 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>92</ID>
<type>AA_AND2</type>
<position>49,-90.5</position>
<input>
<ID>IN_0</ID>99 </input>
<input>
<ID>IN_1</ID>86 </input>
<output>
<ID>OUT</ID>89 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>94</ID>
<type>AE_OR2</type>
<position>57,-87</position>
<input>
<ID>IN_0</ID>88 </input>
<input>
<ID>IN_1</ID>89 </input>
<output>
<ID>OUT</ID>96 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>95</ID>
<type>BE_JKFF_LOW_NT</type>
<position>67.5,-87</position>
<input>
<ID>J</ID>91 </input>
<input>
<ID>K</ID>91 </input>
<output>
<ID>Q</ID>105 </output>
<input>
<ID>clock</ID>96 </input>
<output>
<ID>nQ</ID>93 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>96</ID>
<type>AA_AND2</type>
<position>78.5,-84</position>
<input>
<ID>IN_0</ID>100 </input>
<input>
<ID>IN_1</ID>105 </input>
<output>
<ID>OUT</ID>94 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>97</ID>
<type>AA_AND2</type>
<position>79,-90</position>
<input>
<ID>IN_0</ID>99 </input>
<input>
<ID>IN_1</ID>93 </input>
<output>
<ID>OUT</ID>95 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>98</ID>
<type>AE_OR2</type>
<position>87,-86.5</position>
<input>
<ID>IN_0</ID>94 </input>
<input>
<ID>IN_1</ID>95 </input>
<output>
<ID>OUT</ID>98 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>99</ID>
<type>DA_FROM</type>
<position>61.5,-80.5</position>
<input>
<ID>IN_0</ID>91 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID 1</lparam></gate>
<gate>
<ID>100</ID>
<type>BE_JKFF_LOW_NT</type>
<position>98.5,-86.5</position>
<input>
<ID>J</ID>97 </input>
<input>
<ID>K</ID>97 </input>
<output>
<ID>Q</ID>104 </output>
<input>
<ID>clock</ID>98 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>101</ID>
<type>DA_FROM</type>
<position>92.5,-81</position>
<input>
<ID>IN_0</ID>97 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID 1</lparam></gate>
<gate>
<ID>103</ID>
<type>AA_TOGGLE</type>
<position>26,-75</position>
<output>
<ID>OUT_0</ID>99 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>105</ID>
<type>AE_SMALL_INVERTER</type>
<position>36,-77.5</position>
<input>
<ID>IN_0</ID>99 </input>
<output>
<ID>OUT_0</ID>100 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>114</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>126.5,-68.5</position>
<input>
<ID>IN_0</ID>106 </input>
<input>
<ID>IN_1</ID>105 </input>
<input>
<ID>IN_2</ID>104 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>116</ID>
<type>DE_TO</type>
<position>53.5,-72</position>
<input>
<ID>IN_0</ID>106 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Q1</lparam></gate>
<gate>
<ID>117</ID>
<type>DE_TO</type>
<position>80.5,-72</position>
<input>
<ID>IN_0</ID>105 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Q2</lparam></gate>
<gate>
<ID>118</ID>
<type>DE_TO</type>
<position>107.5,-72</position>
<input>
<ID>IN_0</ID>104 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Q3</lparam></gate>
<gate>
<ID>140</ID>
<type>AE_DFF_LOW_NT</type>
<position>34,-127</position>
<input>
<ID>IN_0</ID>124 </input>
<output>
<ID>OUT_0</ID>125 </output>
<input>
<ID>clear</ID>132 </input>
<input>
<ID>clock</ID>131 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>142</ID>
<type>AE_DFF_LOW_NT</type>
<position>50,-127</position>
<input>
<ID>IN_0</ID>126 </input>
<output>
<ID>OUT_0</ID>127 </output>
<input>
<ID>clear</ID>132 </input>
<input>
<ID>clock</ID>131 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>143</ID>
<type>AE_DFF_LOW_NT</type>
<position>63.5,-127</position>
<input>
<ID>IN_0</ID>128 </input>
<output>
<ID>OUT_0</ID>129 </output>
<input>
<ID>clear</ID>132 </input>
<input>
<ID>clock</ID>131 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>144</ID>
<type>AE_DFF_LOW_NT</type>
<position>79.5,-127</position>
<input>
<ID>IN_0</ID>130 </input>
<output>
<ID>OUTINV_0</ID>124 </output>
<output>
<ID>OUT_0</ID>134 </output>
<input>
<ID>clear</ID>132 </input>
<input>
<ID>clock</ID>131 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>146</ID>
<type>GA_LED</type>
<position>40,-125</position>
<input>
<ID>N_in0</ID>125 </input>
<input>
<ID>N_in1</ID>126 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>149</ID>
<type>GA_LED</type>
<position>57,-125</position>
<input>
<ID>N_in0</ID>127 </input>
<input>
<ID>N_in1</ID>128 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>150</ID>
<type>GA_LED</type>
<position>71.5,-125</position>
<input>
<ID>N_in0</ID>129 </input>
<input>
<ID>N_in1</ID>130 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>151</ID>
<type>BB_CLOCK</type>
<position>22.5,-133.5</position>
<output>
<ID>CLK</ID>131 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>153</ID>
<type>AA_TOGGLE</type>
<position>25,-140.5</position>
<output>
<ID>OUT_0</ID>132 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>154</ID>
<type>GA_LED</type>
<position>85,-125</position>
<input>
<ID>N_in0</ID>134 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>155</ID>
<type>AA_LABEL</type>
<position>35,-111.5</position>
<gparam>LABEL_TEXT 4) Twisted Ring Counter(Jhonson Counter)</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>156</ID>
<type>AA_LABEL</type>
<position>18,-133</position>
<gparam>LABEL_TEXT clock</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>157</ID>
<type>AA_LABEL</type>
<position>21,-140</position>
<gparam>LABEL_TEXT clear</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30,-26,41,-26</points>
<connection>
<GID>4</GID>
<name>CLK</name></connection>
<connection>
<GID>2</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65,-28,65,-23</points>
<connection>
<GID>19</GID>
<name>IN_0</name></connection>
<intersection>-28 2</intersection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>65,-24,67,-24</points>
<connection>
<GID>11</GID>
<name>J</name></connection>
<intersection>65 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>65,-28,67,-28</points>
<connection>
<GID>11</GID>
<name>K</name></connection>
<intersection>65 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15.5,14,22.5,14</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<connection>
<GID>14</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,-28,39,-21.5</points>
<intersection>-28 4</intersection>
<intersection>-24 5</intersection>
<intersection>-21.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>35.5,-21.5,39,-21.5</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>39 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>39,-28,41,-28</points>
<connection>
<GID>2</GID>
<name>K</name></connection>
<intersection>39 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>39,-24,41,-24</points>
<connection>
<GID>2</GID>
<name>J</name></connection>
<intersection>39 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70.5,-21,71.5,-21</points>
<connection>
<GID>25</GID>
<name>N_in0</name></connection>
<intersection>71.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>71.5,-24,71.5,-21</points>
<intersection>-24 4</intersection>
<intersection>-21 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>71.5,-24,73,-24</points>
<connection>
<GID>11</GID>
<name>Q</name></connection>
<intersection>71.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52,-28,52,-23</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>-28 3</intersection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>52,-24,53,-24</points>
<connection>
<GID>10</GID>
<name>J</name></connection>
<intersection>52 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>52,-28,53,-28</points>
<connection>
<GID>10</GID>
<name>K</name></connection>
<intersection>52 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60.5,-23,60.5,-13.5</points>
<connection>
<GID>23</GID>
<name>N_in3</name></connection>
<intersection>-13.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>60.5,-13.5,75.5,-13.5</points>
<connection>
<GID>30</GID>
<name>IN_1</name></connection>
<intersection>60.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>71.5,-20,71.5,-12.5</points>
<connection>
<GID>25</GID>
<name>N_in3</name></connection>
<intersection>-12.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>71.5,-12.5,75.5,-12.5</points>
<connection>
<GID>30</GID>
<name>IN_2</name></connection>
<intersection>71.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>47,-24,48,-24</points>
<connection>
<GID>2</GID>
<name>Q</name></connection>
<connection>
<GID>32</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51.5,-26,51.5,-24</points>
<intersection>-26 1</intersection>
<intersection>-24 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>51.5,-26,53,-26</points>
<connection>
<GID>10</GID>
<name>clock</name></connection>
<intersection>51.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>50,-24,51.5,-24</points>
<connection>
<GID>32</GID>
<name>N_in1</name></connection>
<intersection>51.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49,-23,49,-14.5</points>
<connection>
<GID>32</GID>
<name>N_in3</name></connection>
<intersection>-14.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49,-14.5,75.5,-14.5</points>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<intersection>49 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63.5,-26,63.5,-24</points>
<intersection>-26 1</intersection>
<intersection>-24 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63.5,-26,67,-26</points>
<connection>
<GID>11</GID>
<name>clock</name></connection>
<intersection>63.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>61.5,-24,63.5,-24</points>
<connection>
<GID>23</GID>
<name>N_in1</name></connection>
<intersection>63.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>59,-24,59.5,-24</points>
<connection>
<GID>23</GID>
<name>N_in0</name></connection>
<connection>
<GID>10</GID>
<name>Q</name></connection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>25.5,-55,29,-55</points>
<connection>
<GID>73</GID>
<name>clock</name></connection>
<connection>
<GID>72</GID>
<name>CLK</name></connection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,-57,28.5,-50</points>
<connection>
<GID>74</GID>
<name>IN_0</name></connection>
<intersection>-57 4</intersection>
<intersection>-53 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28.5,-53,29,-53</points>
<connection>
<GID>73</GID>
<name>J</name></connection>
<intersection>28.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>28.5,-57,29,-57</points>
<connection>
<GID>73</GID>
<name>K</name></connection>
<intersection>28.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41.5,-56.5,41.5,-49.5</points>
<connection>
<GID>75</GID>
<name>IN_0</name></connection>
<intersection>-56.5 3</intersection>
<intersection>-52.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>41.5,-52.5,42,-52.5</points>
<connection>
<GID>76</GID>
<name>J</name></connection>
<intersection>41.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>41.5,-56.5,42,-56.5</points>
<connection>
<GID>76</GID>
<name>K</name></connection>
<intersection>41.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,-53,35.5,-46.5</points>
<intersection>-53 2</intersection>
<intersection>-46.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35.5,-46.5,65.5,-46.5</points>
<connection>
<GID>79</GID>
<name>IN_0</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35,-53,35.5,-53</points>
<connection>
<GID>73</GID>
<name>Q</name></connection>
<intersection>35.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-52.5,50.5,-45.5</points>
<intersection>-52.5 2</intersection>
<intersection>-45.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-45.5,65.5,-45.5</points>
<connection>
<GID>79</GID>
<name>IN_1</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48,-52.5,50.5,-52.5</points>
<connection>
<GID>76</GID>
<name>Q</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63.5,-52.5,63.5,-44.5</points>
<intersection>-52.5 2</intersection>
<intersection>-44.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63.5,-44.5,65.5,-44.5</points>
<connection>
<GID>79</GID>
<name>IN_2</name></connection>
<intersection>63.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>61.5,-52.5,63.5,-52.5</points>
<connection>
<GID>78</GID>
<name>Q</name></connection>
<intersection>63.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,-57,38.5,-54.5</points>
<intersection>-57 2</intersection>
<intersection>-54.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38.5,-54.5,42,-54.5</points>
<connection>
<GID>76</GID>
<name>clock</name></connection>
<intersection>38.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35,-57,38.5,-57</points>
<connection>
<GID>73</GID>
<name>nQ</name></connection>
<intersection>38.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51.5,-56.5,51.5,-54.5</points>
<intersection>-56.5 2</intersection>
<intersection>-54.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>51.5,-54.5,55.5,-54.5</points>
<connection>
<GID>78</GID>
<name>clock</name></connection>
<intersection>51.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48,-56.5,51.5,-56.5</points>
<connection>
<GID>76</GID>
<name>nQ</name></connection>
<intersection>51.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55,-52.5,55,-49.5</points>
<connection>
<GID>77</GID>
<name>IN_0</name></connection>
<intersection>-52.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55,-52.5,55.5,-52.5</points>
<connection>
<GID>78</GID>
<name>J</name></connection>
<intersection>55 0</intersection>
<intersection>55.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>55.5,-56.5,55.5,-52.5</points>
<connection>
<GID>78</GID>
<name>K</name></connection>
<intersection>-52.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22,-87.5,34.5,-87.5</points>
<connection>
<GID>81</GID>
<name>CLK</name></connection>
<connection>
<GID>82</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,-89.5,32.5,-82.5</points>
<intersection>-89.5 4</intersection>
<intersection>-85.5 1</intersection>
<intersection>-82.5 6</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32.5,-85.5,34.5,-85.5</points>
<connection>
<GID>82</GID>
<name>J</name></connection>
<intersection>32.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>32.5,-89.5,34.5,-89.5</points>
<connection>
<GID>82</GID>
<name>K</name></connection>
<intersection>32.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>21,-82.5,32.5,-82.5</points>
<connection>
<GID>83</GID>
<name>IN_0</name></connection>
<intersection>32.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43,-91.5,43,-89.5</points>
<intersection>-91.5 1</intersection>
<intersection>-89.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43,-91.5,46,-91.5</points>
<connection>
<GID>92</GID>
<name>IN_1</name></connection>
<intersection>43 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>40.5,-89.5,43,-89.5</points>
<connection>
<GID>82</GID>
<name>nQ</name></connection>
<intersection>43 0</intersection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52.5,-86,52.5,-84.5</points>
<intersection>-86 1</intersection>
<intersection>-84.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>52.5,-86,54,-86</points>
<connection>
<GID>94</GID>
<name>IN_0</name></connection>
<intersection>52.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>51.5,-84.5,52.5,-84.5</points>
<connection>
<GID>91</GID>
<name>OUT</name></connection>
<intersection>52.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53,-90.5,53,-88</points>
<intersection>-90.5 4</intersection>
<intersection>-88 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>53,-88,54,-88</points>
<connection>
<GID>94</GID>
<name>IN_1</name></connection>
<intersection>53 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>52,-90.5,53,-90.5</points>
<connection>
<GID>92</GID>
<name>OUT</name></connection>
<intersection>53 0</intersection></hsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61.5,-89,61.5,-82.5</points>
<connection>
<GID>99</GID>
<name>IN_0</name></connection>
<intersection>-89 4</intersection>
<intersection>-85 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>61.5,-85,64.5,-85</points>
<connection>
<GID>95</GID>
<name>J</name></connection>
<intersection>61.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>61.5,-89,64.5,-89</points>
<connection>
<GID>95</GID>
<name>K</name></connection>
<intersection>61.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,-91,73,-89</points>
<intersection>-91 1</intersection>
<intersection>-89 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73,-91,76,-91</points>
<connection>
<GID>97</GID>
<name>IN_1</name></connection>
<intersection>73 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>70.5,-89,73,-89</points>
<connection>
<GID>95</GID>
<name>nQ</name></connection>
<intersection>73 0</intersection></hsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>82.5,-85.5,82.5,-84</points>
<intersection>-85.5 1</intersection>
<intersection>-84 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>82.5,-85.5,84,-85.5</points>
<connection>
<GID>98</GID>
<name>IN_0</name></connection>
<intersection>82.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>81.5,-84,82.5,-84</points>
<connection>
<GID>96</GID>
<name>OUT</name></connection>
<intersection>82.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83,-90,83,-87.5</points>
<intersection>-90 2</intersection>
<intersection>-87.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>83,-87.5,84,-87.5</points>
<connection>
<GID>98</GID>
<name>IN_1</name></connection>
<intersection>83 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>82,-90,83,-90</points>
<connection>
<GID>97</GID>
<name>OUT</name></connection>
<intersection>83 0</intersection></hsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>60,-87,64.5,-87</points>
<connection>
<GID>95</GID>
<name>clock</name></connection>
<connection>
<GID>94</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>92.5,-88.5,92.5,-83</points>
<connection>
<GID>101</GID>
<name>IN_0</name></connection>
<intersection>-88.5 4</intersection>
<intersection>-84.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>92.5,-84.5,95.5,-84.5</points>
<connection>
<GID>100</GID>
<name>J</name></connection>
<intersection>92.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>92.5,-88.5,95.5,-88.5</points>
<connection>
<GID>100</GID>
<name>K</name></connection>
<intersection>92.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>90,-86.5,95.5,-86.5</points>
<connection>
<GID>100</GID>
<name>clock</name></connection>
<connection>
<GID>98</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28,-75,74,-75</points>
<connection>
<GID>103</GID>
<name>OUT_0</name></connection>
<intersection>32 7</intersection>
<intersection>44 5</intersection>
<intersection>74 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>74,-89,74,-75</points>
<intersection>-89 4</intersection>
<intersection>-75 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>74,-89,76,-89</points>
<connection>
<GID>97</GID>
<name>IN_0</name></connection>
<intersection>74 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>44,-89.5,44,-75</points>
<intersection>-89.5 6</intersection>
<intersection>-75 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>44,-89.5,46,-89.5</points>
<connection>
<GID>92</GID>
<name>IN_0</name></connection>
<intersection>44 5</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>32,-77.5,32,-75</points>
<intersection>-77.5 8</intersection>
<intersection>-75 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>32,-77.5,34,-77.5</points>
<connection>
<GID>105</GID>
<name>IN_0</name></connection>
<intersection>32 7</intersection></hsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38,-77.5,75.5,-77.5</points>
<connection>
<GID>105</GID>
<name>OUT_0</name></connection>
<intersection>45.5 4</intersection>
<intersection>75.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>75.5,-83,75.5,-77.5</points>
<connection>
<GID>96</GID>
<name>IN_0</name></connection>
<intersection>-77.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>45.5,-83.5,45.5,-77.5</points>
<connection>
<GID>91</GID>
<name>IN_0</name></connection>
<intersection>-77.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104,-84.5,104,-67.5</points>
<intersection>-84.5 7</intersection>
<intersection>-72 8</intersection>
<intersection>-67.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>104,-67.5,123.5,-67.5</points>
<connection>
<GID>114</GID>
<name>IN_2</name></connection>
<intersection>104 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>101.5,-84.5,104,-84.5</points>
<connection>
<GID>100</GID>
<name>Q</name></connection>
<intersection>104 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>104,-72,105.5,-72</points>
<connection>
<GID>118</GID>
<name>IN_0</name></connection>
<intersection>104 0</intersection></hsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>75.5,-68.5,123.5,-68.5</points>
<connection>
<GID>114</GID>
<name>IN_1</name></connection>
<intersection>75.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>75.5,-85,75.5,-68.5</points>
<connection>
<GID>96</GID>
<name>IN_1</name></connection>
<intersection>-85 9</intersection>
<intersection>-72 12</intersection>
<intersection>-68.5 6</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>70.5,-85,75.5,-85</points>
<connection>
<GID>95</GID>
<name>Q</name></connection>
<intersection>75.5 8</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>75.5,-72,78.5,-72</points>
<connection>
<GID>117</GID>
<name>IN_0</name></connection>
<intersection>75.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>45.5,-69.5,123.5,-69.5</points>
<connection>
<GID>114</GID>
<name>IN_0</name></connection>
<intersection>45.5 9</intersection>
<intersection>51.5 13</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>45.5,-85.5,45.5,-69.5</points>
<connection>
<GID>91</GID>
<name>IN_1</name></connection>
<intersection>-85.5 10</intersection>
<intersection>-69.5 7</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>40.5,-85.5,45.5,-85.5</points>
<connection>
<GID>82</GID>
<name>Q</name></connection>
<intersection>45.5 9</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>51.5,-72,51.5,-69.5</points>
<connection>
<GID>116</GID>
<name>IN_0</name></connection>
<intersection>-69.5 7</intersection></vsegment></shape></wire>
<wire>
<ID>124</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27,-118,88,-118</points>
<intersection>27 3</intersection>
<intersection>88 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>27,-125,27,-118</points>
<intersection>-125 5</intersection>
<intersection>-118 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>88,-128,88,-118</points>
<intersection>-128 6</intersection>
<intersection>-118 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>27,-125,31,-125</points>
<connection>
<GID>140</GID>
<name>IN_0</name></connection>
<intersection>27 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>82.5,-128,88,-128</points>
<connection>
<GID>144</GID>
<name>OUTINV_0</name></connection>
<intersection>88 4</intersection></hsegment></shape></wire>
<wire>
<ID>125</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>37,-125,39,-125</points>
<connection>
<GID>140</GID>
<name>OUT_0</name></connection>
<connection>
<GID>146</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>126</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41,-125,47,-125</points>
<connection>
<GID>142</GID>
<name>IN_0</name></connection>
<connection>
<GID>146</GID>
<name>N_in1</name></connection></hsegment></shape></wire>
<wire>
<ID>127</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-125,56,-125</points>
<connection>
<GID>142</GID>
<name>OUT_0</name></connection>
<connection>
<GID>149</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>128</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>58,-125,60.5,-125</points>
<connection>
<GID>143</GID>
<name>IN_0</name></connection>
<connection>
<GID>149</GID>
<name>N_in1</name></connection></hsegment></shape></wire>
<wire>
<ID>129</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>66.5,-125,70.5,-125</points>
<connection>
<GID>143</GID>
<name>OUT_0</name></connection>
<connection>
<GID>150</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>130</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>72.5,-125,76.5,-125</points>
<connection>
<GID>144</GID>
<name>IN_0</name></connection>
<connection>
<GID>150</GID>
<name>N_in1</name></connection></hsegment></shape></wire>
<wire>
<ID>131</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-133.5,71.5,-133.5</points>
<connection>
<GID>151</GID>
<name>CLK</name></connection>
<intersection>29 5</intersection>
<intersection>44 4</intersection>
<intersection>57.5 8</intersection>
<intersection>71.5 10</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>44,-133.5,44,-128</points>
<intersection>-133.5 1</intersection>
<intersection>-128 11</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>29,-133.5,29,-128</points>
<intersection>-133.5 1</intersection>
<intersection>-128 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>29,-128,31,-128</points>
<connection>
<GID>140</GID>
<name>clock</name></connection>
<intersection>29 5</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>57.5,-133.5,57.5,-128</points>
<intersection>-133.5 1</intersection>
<intersection>-128 11</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>71.5,-133.5,71.5,-128</points>
<intersection>-133.5 1</intersection>
<intersection>-128 13</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>44,-128,60.5,-128</points>
<connection>
<GID>142</GID>
<name>clock</name></connection>
<connection>
<GID>143</GID>
<name>clock</name></connection>
<intersection>44 4</intersection>
<intersection>57.5 8</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>71.5,-128,76.5,-128</points>
<connection>
<GID>144</GID>
<name>clock</name></connection>
<intersection>71.5 10</intersection></hsegment></shape></wire>
<wire>
<ID>132</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79.5,-140.5,79.5,-131</points>
<connection>
<GID>144</GID>
<name>clear</name></connection>
<intersection>-140.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27,-140.5,79.5,-140.5</points>
<connection>
<GID>153</GID>
<name>OUT_0</name></connection>
<intersection>34 4</intersection>
<intersection>50 3</intersection>
<intersection>63.5 2</intersection>
<intersection>79.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>63.5,-140.5,63.5,-131</points>
<connection>
<GID>143</GID>
<name>clear</name></connection>
<intersection>-140.5 1</intersection></vsegment>
<vsegment>
<ID>3</ID>
<points>50,-140.5,50,-131</points>
<connection>
<GID>142</GID>
<name>clear</name></connection>
<intersection>-140.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>34,-140.5,34,-131</points>
<connection>
<GID>140</GID>
<name>clear</name></connection>
<intersection>-140.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>134</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>82.5,-125,84,-125</points>
<connection>
<GID>144</GID>
<name>OUT_0</name></connection>
<connection>
<GID>154</GID>
<name>N_in0</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 1>
<page 2>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 2>
<page 3>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 3>
<page 4>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 4>
<page 5>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 5>
<page 6>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 6>
<page 7>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 7>
<page 8>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 8>
<page 9>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 9></circuit>